// Verilog netlist created by TD v4.6.116866
// Sun Nov 16 22:07:49 2025

`timescale 1ns / 1ps
module sample_memory  // al_ip/sample_memory.v(14)
  (
  addra,
  addrb,
  cea,
  clka,
  clkb,
  dia,
  dob
  );

  input [12:0] addra;  // al_ip/sample_memory.v(23)
  input [12:0] addrb;  // al_ip/sample_memory.v(24)
  input cea;  // al_ip/sample_memory.v(25)
  input clka;  // al_ip/sample_memory.v(26)
  input clkb;  // al_ip/sample_memory.v(27)
  input [31:0] dia;  // al_ip/sample_memory.v(22)
  output [31:0] dob;  // al_ip/sample_memory.v(19)


  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_000 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,dia[0],open_n14}),
    .dob({open_n39,open_n40,open_n41,open_n42,open_n43,open_n44,open_n45,open_n46,dob[0]}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_001 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n54,open_n55,open_n56,open_n57,open_n58,open_n59,open_n60,dia[1],open_n61}),
    .dob({open_n86,open_n87,open_n88,open_n89,open_n90,open_n91,open_n92,open_n93,dob[1]}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_002 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n101,open_n102,open_n103,open_n104,open_n105,open_n106,open_n107,dia[2],open_n108}),
    .dob({open_n133,open_n134,open_n135,open_n136,open_n137,open_n138,open_n139,open_n140,dob[2]}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_003 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,open_n154,dia[3],open_n155}),
    .dob({open_n180,open_n181,open_n182,open_n183,open_n184,open_n185,open_n186,open_n187,dob[3]}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_004 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n195,open_n196,open_n197,open_n198,open_n199,open_n200,open_n201,dia[4],open_n202}),
    .dob({open_n227,open_n228,open_n229,open_n230,open_n231,open_n232,open_n233,open_n234,dob[4]}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_005 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n242,open_n243,open_n244,open_n245,open_n246,open_n247,open_n248,dia[5],open_n249}),
    .dob({open_n274,open_n275,open_n276,open_n277,open_n278,open_n279,open_n280,open_n281,dob[5]}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_006 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n289,open_n290,open_n291,open_n292,open_n293,open_n294,open_n295,dia[6],open_n296}),
    .dob({open_n321,open_n322,open_n323,open_n324,open_n325,open_n326,open_n327,open_n328,dob[6]}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_007 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n336,open_n337,open_n338,open_n339,open_n340,open_n341,open_n342,dia[7],open_n343}),
    .dob({open_n368,open_n369,open_n370,open_n371,open_n372,open_n373,open_n374,open_n375,dob[7]}));
  // address_offset=0;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_008 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n383,open_n384,open_n385,open_n386,open_n387,open_n388,open_n389,dia[8],open_n390}),
    .dob({open_n415,open_n416,open_n417,open_n418,open_n419,open_n420,open_n421,open_n422,dob[8]}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_009 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n430,open_n431,open_n432,open_n433,open_n434,open_n435,open_n436,dia[9],open_n437}),
    .dob({open_n462,open_n463,open_n464,open_n465,open_n466,open_n467,open_n468,open_n469,dob[9]}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_010 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n477,open_n478,open_n479,open_n480,open_n481,open_n482,open_n483,dia[10],open_n484}),
    .dob({open_n509,open_n510,open_n511,open_n512,open_n513,open_n514,open_n515,open_n516,dob[10]}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_011 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n524,open_n525,open_n526,open_n527,open_n528,open_n529,open_n530,dia[11],open_n531}),
    .dob({open_n556,open_n557,open_n558,open_n559,open_n560,open_n561,open_n562,open_n563,dob[11]}));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_012 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n571,open_n572,open_n573,open_n574,open_n575,open_n576,open_n577,dia[12],open_n578}),
    .dob({open_n603,open_n604,open_n605,open_n606,open_n607,open_n608,open_n609,open_n610,dob[12]}));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_013 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n618,open_n619,open_n620,open_n621,open_n622,open_n623,open_n624,dia[13],open_n625}),
    .dob({open_n650,open_n651,open_n652,open_n653,open_n654,open_n655,open_n656,open_n657,dob[13]}));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_014 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n665,open_n666,open_n667,open_n668,open_n669,open_n670,open_n671,dia[14],open_n672}),
    .dob({open_n697,open_n698,open_n699,open_n700,open_n701,open_n702,open_n703,open_n704,dob[14]}));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_015 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n712,open_n713,open_n714,open_n715,open_n716,open_n717,open_n718,dia[15],open_n719}),
    .dob({open_n744,open_n745,open_n746,open_n747,open_n748,open_n749,open_n750,open_n751,dob[15]}));
  // address_offset=0;data_offset=16;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_016 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n759,open_n760,open_n761,open_n762,open_n763,open_n764,open_n765,dia[16],open_n766}),
    .dob({open_n791,open_n792,open_n793,open_n794,open_n795,open_n796,open_n797,open_n798,dob[16]}));
  // address_offset=0;data_offset=17;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_017 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n806,open_n807,open_n808,open_n809,open_n810,open_n811,open_n812,dia[17],open_n813}),
    .dob({open_n838,open_n839,open_n840,open_n841,open_n842,open_n843,open_n844,open_n845,dob[17]}));
  // address_offset=0;data_offset=18;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_018 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n853,open_n854,open_n855,open_n856,open_n857,open_n858,open_n859,dia[18],open_n860}),
    .dob({open_n885,open_n886,open_n887,open_n888,open_n889,open_n890,open_n891,open_n892,dob[18]}));
  // address_offset=0;data_offset=19;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_019 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n900,open_n901,open_n902,open_n903,open_n904,open_n905,open_n906,dia[19],open_n907}),
    .dob({open_n932,open_n933,open_n934,open_n935,open_n936,open_n937,open_n938,open_n939,dob[19]}));
  // address_offset=0;data_offset=20;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_020 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n947,open_n948,open_n949,open_n950,open_n951,open_n952,open_n953,dia[20],open_n954}),
    .dob({open_n979,open_n980,open_n981,open_n982,open_n983,open_n984,open_n985,open_n986,dob[20]}));
  // address_offset=0;data_offset=21;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_021 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n994,open_n995,open_n996,open_n997,open_n998,open_n999,open_n1000,dia[21],open_n1001}),
    .dob({open_n1026,open_n1027,open_n1028,open_n1029,open_n1030,open_n1031,open_n1032,open_n1033,dob[21]}));
  // address_offset=0;data_offset=22;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_022 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1041,open_n1042,open_n1043,open_n1044,open_n1045,open_n1046,open_n1047,dia[22],open_n1048}),
    .dob({open_n1073,open_n1074,open_n1075,open_n1076,open_n1077,open_n1078,open_n1079,open_n1080,dob[22]}));
  // address_offset=0;data_offset=23;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_023 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1088,open_n1089,open_n1090,open_n1091,open_n1092,open_n1093,open_n1094,dia[23],open_n1095}),
    .dob({open_n1120,open_n1121,open_n1122,open_n1123,open_n1124,open_n1125,open_n1126,open_n1127,dob[23]}));
  // address_offset=0;data_offset=24;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_024 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1135,open_n1136,open_n1137,open_n1138,open_n1139,open_n1140,open_n1141,dia[24],open_n1142}),
    .dob({open_n1167,open_n1168,open_n1169,open_n1170,open_n1171,open_n1172,open_n1173,open_n1174,dob[24]}));
  // address_offset=0;data_offset=25;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_025 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1182,open_n1183,open_n1184,open_n1185,open_n1186,open_n1187,open_n1188,dia[25],open_n1189}),
    .dob({open_n1214,open_n1215,open_n1216,open_n1217,open_n1218,open_n1219,open_n1220,open_n1221,dob[25]}));
  // address_offset=0;data_offset=26;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_026 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1229,open_n1230,open_n1231,open_n1232,open_n1233,open_n1234,open_n1235,dia[26],open_n1236}),
    .dob({open_n1261,open_n1262,open_n1263,open_n1264,open_n1265,open_n1266,open_n1267,open_n1268,dob[26]}));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_027 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1276,open_n1277,open_n1278,open_n1279,open_n1280,open_n1281,open_n1282,dia[27],open_n1283}),
    .dob({open_n1308,open_n1309,open_n1310,open_n1311,open_n1312,open_n1313,open_n1314,open_n1315,dob[27]}));
  // address_offset=0;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_028 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1323,open_n1324,open_n1325,open_n1326,open_n1327,open_n1328,open_n1329,dia[28],open_n1330}),
    .dob({open_n1355,open_n1356,open_n1357,open_n1358,open_n1359,open_n1360,open_n1361,open_n1362,dob[28]}));
  // address_offset=0;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_029 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1370,open_n1371,open_n1372,open_n1373,open_n1374,open_n1375,open_n1376,dia[29],open_n1377}),
    .dob({open_n1402,open_n1403,open_n1404,open_n1405,open_n1406,open_n1407,open_n1408,open_n1409,dob[29]}));
  // address_offset=0;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_030 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1417,open_n1418,open_n1419,open_n1420,open_n1421,open_n1422,open_n1423,dia[30],open_n1424}),
    .dob({open_n1449,open_n1450,open_n1451,open_n1452,open_n1453,open_n1454,open_n1455,open_n1456,dob[30]}));
  // address_offset=0;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_031 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n1464,open_n1465,open_n1466,open_n1467,open_n1468,open_n1469,open_n1470,dia[31],open_n1471}),
    .dob({open_n1496,open_n1497,open_n1498,open_n1499,open_n1500,open_n1501,open_n1502,open_n1503,dob[31]}));

endmodule 

