// Verilog netlist created by TD v4.6.116866
// Wed Nov 19 17:00:13 2025

`timescale 1ns / 1ps
module sample_memory  // al_ip/sample_memory.v(14)
  (
  addra,
  addrb,
  cea,
  clka,
  clkb,
  dia,
  dob
  );

  input [12:0] addra;  // al_ip/sample_memory.v(23)
  input [12:0] addrb;  // al_ip/sample_memory.v(24)
  input cea;  // al_ip/sample_memory.v(25)
  input clka;  // al_ip/sample_memory.v(26)
  input clkb;  // al_ip/sample_memory.v(27)
  input [31:0] dia;  // al_ip/sample_memory.v(22)
  output [31:0] dob;  // al_ip/sample_memory.v(19)

  wire [0:2] addrb_piped;
  wire  \inst_dob_mux_b0/B0_0 ;
  wire  \inst_dob_mux_b0/B0_1 ;
  wire  \inst_dob_mux_b0/B0_2 ;
  wire  \inst_dob_mux_b0/B0_3 ;
  wire  \inst_dob_mux_b0/B1_0 ;
  wire  \inst_dob_mux_b0/B1_1 ;
  wire  \inst_dob_mux_b1/B0_0 ;
  wire  \inst_dob_mux_b1/B0_1 ;
  wire  \inst_dob_mux_b1/B0_2 ;
  wire  \inst_dob_mux_b1/B0_3 ;
  wire  \inst_dob_mux_b1/B1_0 ;
  wire  \inst_dob_mux_b1/B1_1 ;
  wire  \inst_dob_mux_b10/B0_0 ;
  wire  \inst_dob_mux_b10/B0_1 ;
  wire  \inst_dob_mux_b10/B0_2 ;
  wire  \inst_dob_mux_b10/B0_3 ;
  wire  \inst_dob_mux_b10/B1_0 ;
  wire  \inst_dob_mux_b10/B1_1 ;
  wire  \inst_dob_mux_b11/B0_0 ;
  wire  \inst_dob_mux_b11/B0_1 ;
  wire  \inst_dob_mux_b11/B0_2 ;
  wire  \inst_dob_mux_b11/B0_3 ;
  wire  \inst_dob_mux_b11/B1_0 ;
  wire  \inst_dob_mux_b11/B1_1 ;
  wire  \inst_dob_mux_b12/B0_0 ;
  wire  \inst_dob_mux_b12/B0_1 ;
  wire  \inst_dob_mux_b12/B0_2 ;
  wire  \inst_dob_mux_b12/B0_3 ;
  wire  \inst_dob_mux_b12/B1_0 ;
  wire  \inst_dob_mux_b12/B1_1 ;
  wire  \inst_dob_mux_b13/B0_0 ;
  wire  \inst_dob_mux_b13/B0_1 ;
  wire  \inst_dob_mux_b13/B0_2 ;
  wire  \inst_dob_mux_b13/B0_3 ;
  wire  \inst_dob_mux_b13/B1_0 ;
  wire  \inst_dob_mux_b13/B1_1 ;
  wire  \inst_dob_mux_b14/B0_0 ;
  wire  \inst_dob_mux_b14/B0_1 ;
  wire  \inst_dob_mux_b14/B0_2 ;
  wire  \inst_dob_mux_b14/B0_3 ;
  wire  \inst_dob_mux_b14/B1_0 ;
  wire  \inst_dob_mux_b14/B1_1 ;
  wire  \inst_dob_mux_b15/B0_0 ;
  wire  \inst_dob_mux_b15/B0_1 ;
  wire  \inst_dob_mux_b15/B0_2 ;
  wire  \inst_dob_mux_b15/B0_3 ;
  wire  \inst_dob_mux_b15/B1_0 ;
  wire  \inst_dob_mux_b15/B1_1 ;
  wire  \inst_dob_mux_b16/B0_0 ;
  wire  \inst_dob_mux_b16/B0_1 ;
  wire  \inst_dob_mux_b16/B0_2 ;
  wire  \inst_dob_mux_b16/B0_3 ;
  wire  \inst_dob_mux_b16/B1_0 ;
  wire  \inst_dob_mux_b16/B1_1 ;
  wire  \inst_dob_mux_b17/B0_0 ;
  wire  \inst_dob_mux_b17/B0_1 ;
  wire  \inst_dob_mux_b17/B0_2 ;
  wire  \inst_dob_mux_b17/B0_3 ;
  wire  \inst_dob_mux_b17/B1_0 ;
  wire  \inst_dob_mux_b17/B1_1 ;
  wire  \inst_dob_mux_b18/B0_0 ;
  wire  \inst_dob_mux_b18/B0_1 ;
  wire  \inst_dob_mux_b18/B0_2 ;
  wire  \inst_dob_mux_b18/B0_3 ;
  wire  \inst_dob_mux_b18/B1_0 ;
  wire  \inst_dob_mux_b18/B1_1 ;
  wire  \inst_dob_mux_b19/B0_0 ;
  wire  \inst_dob_mux_b19/B0_1 ;
  wire  \inst_dob_mux_b19/B0_2 ;
  wire  \inst_dob_mux_b19/B0_3 ;
  wire  \inst_dob_mux_b19/B1_0 ;
  wire  \inst_dob_mux_b19/B1_1 ;
  wire  \inst_dob_mux_b2/B0_0 ;
  wire  \inst_dob_mux_b2/B0_1 ;
  wire  \inst_dob_mux_b2/B0_2 ;
  wire  \inst_dob_mux_b2/B0_3 ;
  wire  \inst_dob_mux_b2/B1_0 ;
  wire  \inst_dob_mux_b2/B1_1 ;
  wire  \inst_dob_mux_b20/B0_0 ;
  wire  \inst_dob_mux_b20/B0_1 ;
  wire  \inst_dob_mux_b20/B0_2 ;
  wire  \inst_dob_mux_b20/B0_3 ;
  wire  \inst_dob_mux_b20/B1_0 ;
  wire  \inst_dob_mux_b20/B1_1 ;
  wire  \inst_dob_mux_b21/B0_0 ;
  wire  \inst_dob_mux_b21/B0_1 ;
  wire  \inst_dob_mux_b21/B0_2 ;
  wire  \inst_dob_mux_b21/B0_3 ;
  wire  \inst_dob_mux_b21/B1_0 ;
  wire  \inst_dob_mux_b21/B1_1 ;
  wire  \inst_dob_mux_b22/B0_0 ;
  wire  \inst_dob_mux_b22/B0_1 ;
  wire  \inst_dob_mux_b22/B0_2 ;
  wire  \inst_dob_mux_b22/B0_3 ;
  wire  \inst_dob_mux_b22/B1_0 ;
  wire  \inst_dob_mux_b22/B1_1 ;
  wire  \inst_dob_mux_b23/B0_0 ;
  wire  \inst_dob_mux_b23/B0_1 ;
  wire  \inst_dob_mux_b23/B0_2 ;
  wire  \inst_dob_mux_b23/B0_3 ;
  wire  \inst_dob_mux_b23/B1_0 ;
  wire  \inst_dob_mux_b23/B1_1 ;
  wire  \inst_dob_mux_b24/B0_0 ;
  wire  \inst_dob_mux_b24/B0_1 ;
  wire  \inst_dob_mux_b24/B0_2 ;
  wire  \inst_dob_mux_b24/B0_3 ;
  wire  \inst_dob_mux_b24/B1_0 ;
  wire  \inst_dob_mux_b24/B1_1 ;
  wire  \inst_dob_mux_b25/B0_0 ;
  wire  \inst_dob_mux_b25/B0_1 ;
  wire  \inst_dob_mux_b25/B0_2 ;
  wire  \inst_dob_mux_b25/B0_3 ;
  wire  \inst_dob_mux_b25/B1_0 ;
  wire  \inst_dob_mux_b25/B1_1 ;
  wire  \inst_dob_mux_b26/B0_0 ;
  wire  \inst_dob_mux_b26/B0_1 ;
  wire  \inst_dob_mux_b26/B0_2 ;
  wire  \inst_dob_mux_b26/B0_3 ;
  wire  \inst_dob_mux_b26/B1_0 ;
  wire  \inst_dob_mux_b26/B1_1 ;
  wire  \inst_dob_mux_b27/B0_0 ;
  wire  \inst_dob_mux_b27/B0_1 ;
  wire  \inst_dob_mux_b27/B0_2 ;
  wire  \inst_dob_mux_b27/B0_3 ;
  wire  \inst_dob_mux_b27/B1_0 ;
  wire  \inst_dob_mux_b27/B1_1 ;
  wire  \inst_dob_mux_b28/B0_0 ;
  wire  \inst_dob_mux_b28/B0_1 ;
  wire  \inst_dob_mux_b28/B0_2 ;
  wire  \inst_dob_mux_b28/B0_3 ;
  wire  \inst_dob_mux_b28/B1_0 ;
  wire  \inst_dob_mux_b28/B1_1 ;
  wire  \inst_dob_mux_b29/B0_0 ;
  wire  \inst_dob_mux_b29/B0_1 ;
  wire  \inst_dob_mux_b29/B0_2 ;
  wire  \inst_dob_mux_b29/B0_3 ;
  wire  \inst_dob_mux_b29/B1_0 ;
  wire  \inst_dob_mux_b29/B1_1 ;
  wire  \inst_dob_mux_b3/B0_0 ;
  wire  \inst_dob_mux_b3/B0_1 ;
  wire  \inst_dob_mux_b3/B0_2 ;
  wire  \inst_dob_mux_b3/B0_3 ;
  wire  \inst_dob_mux_b3/B1_0 ;
  wire  \inst_dob_mux_b3/B1_1 ;
  wire  \inst_dob_mux_b30/B0_0 ;
  wire  \inst_dob_mux_b30/B0_1 ;
  wire  \inst_dob_mux_b30/B0_2 ;
  wire  \inst_dob_mux_b30/B0_3 ;
  wire  \inst_dob_mux_b30/B1_0 ;
  wire  \inst_dob_mux_b30/B1_1 ;
  wire  \inst_dob_mux_b31/B0_0 ;
  wire  \inst_dob_mux_b31/B0_1 ;
  wire  \inst_dob_mux_b31/B0_2 ;
  wire  \inst_dob_mux_b31/B0_3 ;
  wire  \inst_dob_mux_b31/B1_0 ;
  wire  \inst_dob_mux_b31/B1_1 ;
  wire  \inst_dob_mux_b4/B0_0 ;
  wire  \inst_dob_mux_b4/B0_1 ;
  wire  \inst_dob_mux_b4/B0_2 ;
  wire  \inst_dob_mux_b4/B0_3 ;
  wire  \inst_dob_mux_b4/B1_0 ;
  wire  \inst_dob_mux_b4/B1_1 ;
  wire  \inst_dob_mux_b5/B0_0 ;
  wire  \inst_dob_mux_b5/B0_1 ;
  wire  \inst_dob_mux_b5/B0_2 ;
  wire  \inst_dob_mux_b5/B0_3 ;
  wire  \inst_dob_mux_b5/B1_0 ;
  wire  \inst_dob_mux_b5/B1_1 ;
  wire  \inst_dob_mux_b6/B0_0 ;
  wire  \inst_dob_mux_b6/B0_1 ;
  wire  \inst_dob_mux_b6/B0_2 ;
  wire  \inst_dob_mux_b6/B0_3 ;
  wire  \inst_dob_mux_b6/B1_0 ;
  wire  \inst_dob_mux_b6/B1_1 ;
  wire  \inst_dob_mux_b7/B0_0 ;
  wire  \inst_dob_mux_b7/B0_1 ;
  wire  \inst_dob_mux_b7/B0_2 ;
  wire  \inst_dob_mux_b7/B0_3 ;
  wire  \inst_dob_mux_b7/B1_0 ;
  wire  \inst_dob_mux_b7/B1_1 ;
  wire  \inst_dob_mux_b8/B0_0 ;
  wire  \inst_dob_mux_b8/B0_1 ;
  wire  \inst_dob_mux_b8/B0_2 ;
  wire  \inst_dob_mux_b8/B0_3 ;
  wire  \inst_dob_mux_b8/B1_0 ;
  wire  \inst_dob_mux_b8/B1_1 ;
  wire  \inst_dob_mux_b9/B0_0 ;
  wire  \inst_dob_mux_b9/B0_1 ;
  wire  \inst_dob_mux_b9/B0_2 ;
  wire  \inst_dob_mux_b9/B0_3 ;
  wire  \inst_dob_mux_b9/B1_0 ;
  wire  \inst_dob_mux_b9/B1_1 ;
  wire inst_dob_i0_000;
  wire inst_dob_i0_001;
  wire inst_dob_i0_002;
  wire inst_dob_i0_003;
  wire inst_dob_i0_004;
  wire inst_dob_i0_005;
  wire inst_dob_i0_006;
  wire inst_dob_i0_007;
  wire inst_dob_i0_008;
  wire inst_dob_i0_009;
  wire inst_dob_i0_010;
  wire inst_dob_i0_011;
  wire inst_dob_i0_012;
  wire inst_dob_i0_013;
  wire inst_dob_i0_014;
  wire inst_dob_i0_015;
  wire inst_dob_i0_016;
  wire inst_dob_i0_017;
  wire inst_dob_i0_018;
  wire inst_dob_i0_019;
  wire inst_dob_i0_020;
  wire inst_dob_i0_021;
  wire inst_dob_i0_022;
  wire inst_dob_i0_023;
  wire inst_dob_i0_024;
  wire inst_dob_i0_025;
  wire inst_dob_i0_026;
  wire inst_dob_i0_027;
  wire inst_dob_i0_028;
  wire inst_dob_i0_029;
  wire inst_dob_i0_030;
  wire inst_dob_i0_031;
  wire inst_dob_i1_000;
  wire inst_dob_i1_001;
  wire inst_dob_i1_002;
  wire inst_dob_i1_003;
  wire inst_dob_i1_004;
  wire inst_dob_i1_005;
  wire inst_dob_i1_006;
  wire inst_dob_i1_007;
  wire inst_dob_i1_008;
  wire inst_dob_i1_009;
  wire inst_dob_i1_010;
  wire inst_dob_i1_011;
  wire inst_dob_i1_012;
  wire inst_dob_i1_013;
  wire inst_dob_i1_014;
  wire inst_dob_i1_015;
  wire inst_dob_i1_016;
  wire inst_dob_i1_017;
  wire inst_dob_i1_018;
  wire inst_dob_i1_019;
  wire inst_dob_i1_020;
  wire inst_dob_i1_021;
  wire inst_dob_i1_022;
  wire inst_dob_i1_023;
  wire inst_dob_i1_024;
  wire inst_dob_i1_025;
  wire inst_dob_i1_026;
  wire inst_dob_i2_000;
  wire inst_dob_i2_001;
  wire inst_dob_i2_002;
  wire inst_dob_i2_003;
  wire inst_dob_i2_004;
  wire inst_dob_i2_005;
  wire inst_dob_i2_006;
  wire inst_dob_i2_007;
  wire inst_dob_i2_008;
  wire inst_dob_i2_009;
  wire inst_dob_i2_010;
  wire inst_dob_i2_011;
  wire inst_dob_i2_012;
  wire inst_dob_i2_013;
  wire inst_dob_i2_014;
  wire inst_dob_i2_015;
  wire inst_dob_i2_016;
  wire inst_dob_i2_017;
  wire inst_dob_i2_018;
  wire inst_dob_i2_019;
  wire inst_dob_i2_020;
  wire inst_dob_i2_021;
  wire inst_dob_i2_022;
  wire inst_dob_i2_023;
  wire inst_dob_i2_024;
  wire inst_dob_i2_025;
  wire inst_dob_i2_026;
  wire inst_dob_i3_000;
  wire inst_dob_i3_001;
  wire inst_dob_i3_002;
  wire inst_dob_i3_003;
  wire inst_dob_i3_004;
  wire inst_dob_i3_005;
  wire inst_dob_i3_006;
  wire inst_dob_i3_007;
  wire inst_dob_i3_008;
  wire inst_dob_i3_009;
  wire inst_dob_i3_010;
  wire inst_dob_i3_011;
  wire inst_dob_i3_012;
  wire inst_dob_i3_013;
  wire inst_dob_i3_014;
  wire inst_dob_i3_015;
  wire inst_dob_i3_016;
  wire inst_dob_i3_017;
  wire inst_dob_i3_018;
  wire inst_dob_i3_019;
  wire inst_dob_i3_020;
  wire inst_dob_i3_021;
  wire inst_dob_i3_022;
  wire inst_dob_i3_023;
  wire inst_dob_i3_024;
  wire inst_dob_i3_025;
  wire inst_dob_i3_026;
  wire inst_dob_i4_000;
  wire inst_dob_i4_001;
  wire inst_dob_i4_002;
  wire inst_dob_i4_003;
  wire inst_dob_i4_004;
  wire inst_dob_i4_005;
  wire inst_dob_i4_006;
  wire inst_dob_i4_007;
  wire inst_dob_i4_008;
  wire inst_dob_i4_009;
  wire inst_dob_i4_010;
  wire inst_dob_i4_011;
  wire inst_dob_i4_012;
  wire inst_dob_i4_013;
  wire inst_dob_i4_014;
  wire inst_dob_i4_015;
  wire inst_dob_i4_016;
  wire inst_dob_i4_017;
  wire inst_dob_i4_018;
  wire inst_dob_i4_019;
  wire inst_dob_i4_020;
  wire inst_dob_i4_021;
  wire inst_dob_i4_022;
  wire inst_dob_i4_023;
  wire inst_dob_i4_024;
  wire inst_dob_i4_025;
  wire inst_dob_i4_026;
  wire inst_dob_i5_000;
  wire inst_dob_i5_001;
  wire inst_dob_i5_002;
  wire inst_dob_i5_003;
  wire inst_dob_i5_004;
  wire inst_dob_i5_005;
  wire inst_dob_i5_006;
  wire inst_dob_i5_007;
  wire inst_dob_i5_008;
  wire inst_dob_i5_009;
  wire inst_dob_i5_010;
  wire inst_dob_i5_011;
  wire inst_dob_i5_012;
  wire inst_dob_i5_013;
  wire inst_dob_i5_014;
  wire inst_dob_i5_015;
  wire inst_dob_i5_016;
  wire inst_dob_i5_017;
  wire inst_dob_i5_018;
  wire inst_dob_i5_019;
  wire inst_dob_i5_020;
  wire inst_dob_i5_021;
  wire inst_dob_i5_022;
  wire inst_dob_i5_023;
  wire inst_dob_i5_024;
  wire inst_dob_i5_025;
  wire inst_dob_i5_026;
  wire inst_dob_i6_000;
  wire inst_dob_i6_001;
  wire inst_dob_i6_002;
  wire inst_dob_i6_003;
  wire inst_dob_i6_004;
  wire inst_dob_i6_005;
  wire inst_dob_i6_006;
  wire inst_dob_i6_007;
  wire inst_dob_i6_008;
  wire inst_dob_i6_009;
  wire inst_dob_i6_010;
  wire inst_dob_i6_011;
  wire inst_dob_i6_012;
  wire inst_dob_i6_013;
  wire inst_dob_i6_014;
  wire inst_dob_i6_015;
  wire inst_dob_i6_016;
  wire inst_dob_i6_017;
  wire inst_dob_i6_018;
  wire inst_dob_i6_019;
  wire inst_dob_i6_020;
  wire inst_dob_i6_021;
  wire inst_dob_i6_022;
  wire inst_dob_i6_023;
  wire inst_dob_i6_024;
  wire inst_dob_i6_025;
  wire inst_dob_i6_026;
  wire inst_dob_i7_000;
  wire inst_dob_i7_001;
  wire inst_dob_i7_002;
  wire inst_dob_i7_003;
  wire inst_dob_i7_004;
  wire inst_dob_i7_005;
  wire inst_dob_i7_006;
  wire inst_dob_i7_007;
  wire inst_dob_i7_008;
  wire inst_dob_i7_009;
  wire inst_dob_i7_010;
  wire inst_dob_i7_011;
  wire inst_dob_i7_012;
  wire inst_dob_i7_013;
  wire inst_dob_i7_014;
  wire inst_dob_i7_015;
  wire inst_dob_i7_016;
  wire inst_dob_i7_017;
  wire inst_dob_i7_018;
  wire inst_dob_i7_019;
  wire inst_dob_i7_020;
  wire inst_dob_i7_021;
  wire inst_dob_i7_022;
  wire inst_dob_i7_023;
  wire inst_dob_i7_024;
  wire inst_dob_i7_025;
  wire inst_dob_i7_026;

  reg_ar_as_w1 addrb_pipe_b0 (
    .clk(clkb),
    .d(addrb[10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(addrb_piped[0]));
  reg_ar_as_w1 addrb_pipe_b1 (
    .clk(clkb),
    .d(addrb[11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(addrb_piped[1]));
  reg_ar_as_w1 addrb_pipe_b2 (
    .clk(clkb),
    .d(addrb[12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(addrb_piped[2]));
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i0_008,inst_dob_i0_007,inst_dob_i0_006,inst_dob_i0_005,inst_dob_i0_004,inst_dob_i0_003,inst_dob_i0_002,inst_dob_i0_001,inst_dob_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i0_017,inst_dob_i0_016,inst_dob_i0_015,inst_dob_i0_014,inst_dob_i0_013,inst_dob_i0_012,inst_dob_i0_011,inst_dob_i0_010,inst_dob_i0_009}));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i0_026,inst_dob_i0_025,inst_dob_i0_024,inst_dob_i0_023,inst_dob_i0_022,inst_dob_i0_021,inst_dob_i0_020,inst_dob_i0_019,inst_dob_i0_018}));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_027 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,open_n88,dia[27],open_n89}),
    .dob({open_n114,open_n115,open_n116,open_n117,open_n118,open_n119,open_n120,open_n121,inst_dob_i0_027}));
  // address_offset=0;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_028 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n129,open_n130,open_n131,open_n132,open_n133,open_n134,open_n135,dia[28],open_n136}),
    .dob({open_n161,open_n162,open_n163,open_n164,open_n165,open_n166,open_n167,open_n168,inst_dob_i0_028}));
  // address_offset=0;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_029 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n176,open_n177,open_n178,open_n179,open_n180,open_n181,open_n182,dia[29],open_n183}),
    .dob({open_n208,open_n209,open_n210,open_n211,open_n212,open_n213,open_n214,open_n215,inst_dob_i0_029}));
  // address_offset=0;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_030 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n223,open_n224,open_n225,open_n226,open_n227,open_n228,open_n229,dia[30],open_n230}),
    .dob({open_n255,open_n256,open_n257,open_n258,open_n259,open_n260,open_n261,open_n262,inst_dob_i0_030}));
  // address_offset=0;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_031 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n270,open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,dia[31],open_n277}),
    .dob({open_n302,open_n303,open_n304,open_n305,open_n306,open_n307,open_n308,open_n309,inst_dob_i0_031}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i1_008,inst_dob_i1_007,inst_dob_i1_006,inst_dob_i1_005,inst_dob_i1_004,inst_dob_i1_003,inst_dob_i1_002,inst_dob_i1_001,inst_dob_i1_000}));
  // address_offset=1024;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i1_017,inst_dob_i1_016,inst_dob_i1_015,inst_dob_i1_014,inst_dob_i1_013,inst_dob_i1_012,inst_dob_i1_011,inst_dob_i1_010,inst_dob_i1_009}));
  // address_offset=1024;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i1_026,inst_dob_i1_025,inst_dob_i1_024,inst_dob_i1_023,inst_dob_i1_022,inst_dob_i1_021,inst_dob_i1_020,inst_dob_i1_019,inst_dob_i1_018}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i2_008,inst_dob_i2_007,inst_dob_i2_006,inst_dob_i2_005,inst_dob_i2_004,inst_dob_i2_003,inst_dob_i2_002,inst_dob_i2_001,inst_dob_i2_000}));
  // address_offset=2048;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i2_017,inst_dob_i2_016,inst_dob_i2_015,inst_dob_i2_014,inst_dob_i2_013,inst_dob_i2_012,inst_dob_i2_011,inst_dob_i2_010,inst_dob_i2_009}));
  // address_offset=2048;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i2_026,inst_dob_i2_025,inst_dob_i2_024,inst_dob_i2_023,inst_dob_i2_022,inst_dob_i2_021,inst_dob_i2_020,inst_dob_i2_019,inst_dob_i2_018}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i3_008,inst_dob_i3_007,inst_dob_i3_006,inst_dob_i3_005,inst_dob_i3_004,inst_dob_i3_003,inst_dob_i3_002,inst_dob_i3_001,inst_dob_i3_000}));
  // address_offset=3072;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i3_017,inst_dob_i3_016,inst_dob_i3_015,inst_dob_i3_014,inst_dob_i3_013,inst_dob_i3_012,inst_dob_i3_011,inst_dob_i3_010,inst_dob_i3_009}));
  // address_offset=3072;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i3_026,inst_dob_i3_025,inst_dob_i3_024,inst_dob_i3_023,inst_dob_i3_022,inst_dob_i3_021,inst_dob_i3_020,inst_dob_i3_019,inst_dob_i3_018}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i4_008,inst_dob_i4_007,inst_dob_i4_006,inst_dob_i4_005,inst_dob_i4_004,inst_dob_i4_003,inst_dob_i4_002,inst_dob_i4_001,inst_dob_i4_000}));
  // address_offset=4096;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i4_017,inst_dob_i4_016,inst_dob_i4_015,inst_dob_i4_014,inst_dob_i4_013,inst_dob_i4_012,inst_dob_i4_011,inst_dob_i4_010,inst_dob_i4_009}));
  // address_offset=4096;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i4_026,inst_dob_i4_025,inst_dob_i4_024,inst_dob_i4_023,inst_dob_i4_022,inst_dob_i4_021,inst_dob_i4_020,inst_dob_i4_019,inst_dob_i4_018}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i5_008,inst_dob_i5_007,inst_dob_i5_006,inst_dob_i5_005,inst_dob_i5_004,inst_dob_i5_003,inst_dob_i5_002,inst_dob_i5_001,inst_dob_i5_000}));
  // address_offset=5120;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i5_017,inst_dob_i5_016,inst_dob_i5_015,inst_dob_i5_014,inst_dob_i5_013,inst_dob_i5_012,inst_dob_i5_011,inst_dob_i5_010,inst_dob_i5_009}));
  // address_offset=5120;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i5_026,inst_dob_i5_025,inst_dob_i5_024,inst_dob_i5_023,inst_dob_i5_022,inst_dob_i5_021,inst_dob_i5_020,inst_dob_i5_019,inst_dob_i5_018}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i6_008,inst_dob_i6_007,inst_dob_i6_006,inst_dob_i6_005,inst_dob_i6_004,inst_dob_i6_003,inst_dob_i6_002,inst_dob_i6_001,inst_dob_i6_000}));
  // address_offset=6144;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_006144_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i6_017,inst_dob_i6_016,inst_dob_i6_015,inst_dob_i6_014,inst_dob_i6_013,inst_dob_i6_012,inst_dob_i6_011,inst_dob_i6_010,inst_dob_i6_009}));
  // address_offset=6144;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_006144_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i6_026,inst_dob_i6_025,inst_dob_i6_024,inst_dob_i6_023,inst_dob_i6_022,inst_dob_i6_021,inst_dob_i6_020,inst_dob_i6_019,inst_dob_i6_018}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i7_008,inst_dob_i7_007,inst_dob_i7_006,inst_dob_i7_005,inst_dob_i7_004,inst_dob_i7_003,inst_dob_i7_002,inst_dob_i7_001,inst_dob_i7_000}));
  // address_offset=7168;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_007168_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i7_017,inst_dob_i7_016,inst_dob_i7_015,inst_dob_i7_014,inst_dob_i7_013,inst_dob_i7_012,inst_dob_i7_011,inst_dob_i7_010,inst_dob_i7_009}));
  // address_offset=7168;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_007168_018 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[26:18]),
    .dob({inst_dob_i7_026,inst_dob_i7_025,inst_dob_i7_024,inst_dob_i7_023,inst_dob_i7_022,inst_dob_i7_021,inst_dob_i7_020,inst_dob_i7_019,inst_dob_i7_018}));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_0  (
    .i0(inst_dob_i0_000),
    .i1(inst_dob_i1_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_1  (
    .i0(inst_dob_i2_000),
    .i1(inst_dob_i3_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_2  (
    .i0(inst_dob_i4_000),
    .i1(inst_dob_i5_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_3  (
    .i0(inst_dob_i6_000),
    .i1(inst_dob_i7_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b0/B0_0 ),
    .i1(\inst_dob_mux_b0/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b0/B0_2 ),
    .i1(\inst_dob_mux_b0/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b0/B1_0 ),
    .i1(\inst_dob_mux_b0/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[0]));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_0  (
    .i0(inst_dob_i0_001),
    .i1(inst_dob_i1_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_1  (
    .i0(inst_dob_i2_001),
    .i1(inst_dob_i3_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_2  (
    .i0(inst_dob_i4_001),
    .i1(inst_dob_i5_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_3  (
    .i0(inst_dob_i6_001),
    .i1(inst_dob_i7_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b1/B0_0 ),
    .i1(\inst_dob_mux_b1/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b1/B0_2 ),
    .i1(\inst_dob_mux_b1/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b1/B1_0 ),
    .i1(\inst_dob_mux_b1/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[1]));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_0  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i1_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_1  (
    .i0(inst_dob_i2_010),
    .i1(inst_dob_i3_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_2  (
    .i0(inst_dob_i4_010),
    .i1(inst_dob_i5_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_3  (
    .i0(inst_dob_i6_010),
    .i1(inst_dob_i7_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b10/B0_0 ),
    .i1(\inst_dob_mux_b10/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b10/B0_2 ),
    .i1(\inst_dob_mux_b10/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b10/B1_0 ),
    .i1(\inst_dob_mux_b10/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[10]));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_0  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i1_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_1  (
    .i0(inst_dob_i2_011),
    .i1(inst_dob_i3_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_2  (
    .i0(inst_dob_i4_011),
    .i1(inst_dob_i5_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_3  (
    .i0(inst_dob_i6_011),
    .i1(inst_dob_i7_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b11/B0_0 ),
    .i1(\inst_dob_mux_b11/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b11/B0_2 ),
    .i1(\inst_dob_mux_b11/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b11/B1_0 ),
    .i1(\inst_dob_mux_b11/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[11]));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_0  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i1_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_1  (
    .i0(inst_dob_i2_012),
    .i1(inst_dob_i3_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_2  (
    .i0(inst_dob_i4_012),
    .i1(inst_dob_i5_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_3  (
    .i0(inst_dob_i6_012),
    .i1(inst_dob_i7_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b12/B0_0 ),
    .i1(\inst_dob_mux_b12/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b12/B0_2 ),
    .i1(\inst_dob_mux_b12/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b12/B1_0 ),
    .i1(\inst_dob_mux_b12/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[12]));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_0  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i1_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_1  (
    .i0(inst_dob_i2_013),
    .i1(inst_dob_i3_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_2  (
    .i0(inst_dob_i4_013),
    .i1(inst_dob_i5_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_3  (
    .i0(inst_dob_i6_013),
    .i1(inst_dob_i7_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b13/B0_0 ),
    .i1(\inst_dob_mux_b13/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b13/B0_2 ),
    .i1(\inst_dob_mux_b13/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b13/B1_0 ),
    .i1(\inst_dob_mux_b13/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[13]));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_0  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i1_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_1  (
    .i0(inst_dob_i2_014),
    .i1(inst_dob_i3_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_2  (
    .i0(inst_dob_i4_014),
    .i1(inst_dob_i5_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_3  (
    .i0(inst_dob_i6_014),
    .i1(inst_dob_i7_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b14/B0_0 ),
    .i1(\inst_dob_mux_b14/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b14/B0_2 ),
    .i1(\inst_dob_mux_b14/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b14/B1_0 ),
    .i1(\inst_dob_mux_b14/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[14]));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_0  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i1_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_1  (
    .i0(inst_dob_i2_015),
    .i1(inst_dob_i3_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_2  (
    .i0(inst_dob_i4_015),
    .i1(inst_dob_i5_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_3  (
    .i0(inst_dob_i6_015),
    .i1(inst_dob_i7_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b15/B0_0 ),
    .i1(\inst_dob_mux_b15/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b15/B0_2 ),
    .i1(\inst_dob_mux_b15/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b15/B1_0 ),
    .i1(\inst_dob_mux_b15/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[15]));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_0  (
    .i0(inst_dob_i0_016),
    .i1(inst_dob_i1_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_0 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_1  (
    .i0(inst_dob_i2_016),
    .i1(inst_dob_i3_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_1 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_2  (
    .i0(inst_dob_i4_016),
    .i1(inst_dob_i5_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_2 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_3  (
    .i0(inst_dob_i6_016),
    .i1(inst_dob_i7_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_3 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b16/B0_0 ),
    .i1(\inst_dob_mux_b16/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b16/B1_0 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b16/B0_2 ),
    .i1(\inst_dob_mux_b16/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b16/B1_1 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b16/B1_0 ),
    .i1(\inst_dob_mux_b16/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[16]));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_0  (
    .i0(inst_dob_i0_017),
    .i1(inst_dob_i1_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_0 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_1  (
    .i0(inst_dob_i2_017),
    .i1(inst_dob_i3_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_1 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_2  (
    .i0(inst_dob_i4_017),
    .i1(inst_dob_i5_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_2 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_3  (
    .i0(inst_dob_i6_017),
    .i1(inst_dob_i7_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_3 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b17/B0_0 ),
    .i1(\inst_dob_mux_b17/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b17/B1_0 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b17/B0_2 ),
    .i1(\inst_dob_mux_b17/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b17/B1_1 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b17/B1_0 ),
    .i1(\inst_dob_mux_b17/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[17]));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_0_0  (
    .i0(inst_dob_i0_018),
    .i1(inst_dob_i1_018),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b18/B0_0 ));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_0_1  (
    .i0(inst_dob_i2_018),
    .i1(inst_dob_i3_018),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b18/B0_1 ));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_0_2  (
    .i0(inst_dob_i4_018),
    .i1(inst_dob_i5_018),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b18/B0_2 ));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_0_3  (
    .i0(inst_dob_i6_018),
    .i1(inst_dob_i7_018),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b18/B0_3 ));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b18/B0_0 ),
    .i1(\inst_dob_mux_b18/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b18/B1_0 ));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b18/B0_2 ),
    .i1(\inst_dob_mux_b18/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b18/B1_1 ));
  AL_MUX \inst_dob_mux_b18/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b18/B1_0 ),
    .i1(\inst_dob_mux_b18/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[18]));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_0_0  (
    .i0(inst_dob_i0_019),
    .i1(inst_dob_i1_019),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b19/B0_0 ));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_0_1  (
    .i0(inst_dob_i2_019),
    .i1(inst_dob_i3_019),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b19/B0_1 ));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_0_2  (
    .i0(inst_dob_i4_019),
    .i1(inst_dob_i5_019),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b19/B0_2 ));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_0_3  (
    .i0(inst_dob_i6_019),
    .i1(inst_dob_i7_019),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b19/B0_3 ));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b19/B0_0 ),
    .i1(\inst_dob_mux_b19/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b19/B1_0 ));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b19/B0_2 ),
    .i1(\inst_dob_mux_b19/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b19/B1_1 ));
  AL_MUX \inst_dob_mux_b19/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b19/B1_0 ),
    .i1(\inst_dob_mux_b19/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[19]));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_0  (
    .i0(inst_dob_i0_002),
    .i1(inst_dob_i1_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_1  (
    .i0(inst_dob_i2_002),
    .i1(inst_dob_i3_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_2  (
    .i0(inst_dob_i4_002),
    .i1(inst_dob_i5_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_3  (
    .i0(inst_dob_i6_002),
    .i1(inst_dob_i7_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b2/B0_0 ),
    .i1(\inst_dob_mux_b2/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b2/B0_2 ),
    .i1(\inst_dob_mux_b2/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b2/B1_0 ),
    .i1(\inst_dob_mux_b2/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[2]));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_0_0  (
    .i0(inst_dob_i0_020),
    .i1(inst_dob_i1_020),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b20/B0_0 ));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_0_1  (
    .i0(inst_dob_i2_020),
    .i1(inst_dob_i3_020),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b20/B0_1 ));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_0_2  (
    .i0(inst_dob_i4_020),
    .i1(inst_dob_i5_020),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b20/B0_2 ));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_0_3  (
    .i0(inst_dob_i6_020),
    .i1(inst_dob_i7_020),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b20/B0_3 ));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b20/B0_0 ),
    .i1(\inst_dob_mux_b20/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b20/B1_0 ));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b20/B0_2 ),
    .i1(\inst_dob_mux_b20/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b20/B1_1 ));
  AL_MUX \inst_dob_mux_b20/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b20/B1_0 ),
    .i1(\inst_dob_mux_b20/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[20]));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_0_0  (
    .i0(inst_dob_i0_021),
    .i1(inst_dob_i1_021),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b21/B0_0 ));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_0_1  (
    .i0(inst_dob_i2_021),
    .i1(inst_dob_i3_021),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b21/B0_1 ));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_0_2  (
    .i0(inst_dob_i4_021),
    .i1(inst_dob_i5_021),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b21/B0_2 ));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_0_3  (
    .i0(inst_dob_i6_021),
    .i1(inst_dob_i7_021),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b21/B0_3 ));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b21/B0_0 ),
    .i1(\inst_dob_mux_b21/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b21/B1_0 ));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b21/B0_2 ),
    .i1(\inst_dob_mux_b21/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b21/B1_1 ));
  AL_MUX \inst_dob_mux_b21/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b21/B1_0 ),
    .i1(\inst_dob_mux_b21/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[21]));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_0_0  (
    .i0(inst_dob_i0_022),
    .i1(inst_dob_i1_022),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b22/B0_0 ));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_0_1  (
    .i0(inst_dob_i2_022),
    .i1(inst_dob_i3_022),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b22/B0_1 ));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_0_2  (
    .i0(inst_dob_i4_022),
    .i1(inst_dob_i5_022),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b22/B0_2 ));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_0_3  (
    .i0(inst_dob_i6_022),
    .i1(inst_dob_i7_022),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b22/B0_3 ));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b22/B0_0 ),
    .i1(\inst_dob_mux_b22/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b22/B1_0 ));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b22/B0_2 ),
    .i1(\inst_dob_mux_b22/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b22/B1_1 ));
  AL_MUX \inst_dob_mux_b22/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b22/B1_0 ),
    .i1(\inst_dob_mux_b22/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[22]));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_0_0  (
    .i0(inst_dob_i0_023),
    .i1(inst_dob_i1_023),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b23/B0_0 ));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_0_1  (
    .i0(inst_dob_i2_023),
    .i1(inst_dob_i3_023),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b23/B0_1 ));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_0_2  (
    .i0(inst_dob_i4_023),
    .i1(inst_dob_i5_023),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b23/B0_2 ));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_0_3  (
    .i0(inst_dob_i6_023),
    .i1(inst_dob_i7_023),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b23/B0_3 ));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b23/B0_0 ),
    .i1(\inst_dob_mux_b23/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b23/B1_0 ));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b23/B0_2 ),
    .i1(\inst_dob_mux_b23/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b23/B1_1 ));
  AL_MUX \inst_dob_mux_b23/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b23/B1_0 ),
    .i1(\inst_dob_mux_b23/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[23]));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_0_0  (
    .i0(inst_dob_i0_024),
    .i1(inst_dob_i1_024),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b24/B0_0 ));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_0_1  (
    .i0(inst_dob_i2_024),
    .i1(inst_dob_i3_024),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b24/B0_1 ));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_0_2  (
    .i0(inst_dob_i4_024),
    .i1(inst_dob_i5_024),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b24/B0_2 ));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_0_3  (
    .i0(inst_dob_i6_024),
    .i1(inst_dob_i7_024),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b24/B0_3 ));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b24/B0_0 ),
    .i1(\inst_dob_mux_b24/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b24/B1_0 ));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b24/B0_2 ),
    .i1(\inst_dob_mux_b24/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b24/B1_1 ));
  AL_MUX \inst_dob_mux_b24/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b24/B1_0 ),
    .i1(\inst_dob_mux_b24/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[24]));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_0_0  (
    .i0(inst_dob_i0_025),
    .i1(inst_dob_i1_025),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b25/B0_0 ));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_0_1  (
    .i0(inst_dob_i2_025),
    .i1(inst_dob_i3_025),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b25/B0_1 ));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_0_2  (
    .i0(inst_dob_i4_025),
    .i1(inst_dob_i5_025),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b25/B0_2 ));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_0_3  (
    .i0(inst_dob_i6_025),
    .i1(inst_dob_i7_025),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b25/B0_3 ));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b25/B0_0 ),
    .i1(\inst_dob_mux_b25/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b25/B1_0 ));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b25/B0_2 ),
    .i1(\inst_dob_mux_b25/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b25/B1_1 ));
  AL_MUX \inst_dob_mux_b25/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b25/B1_0 ),
    .i1(\inst_dob_mux_b25/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[25]));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_0_0  (
    .i0(inst_dob_i0_026),
    .i1(inst_dob_i1_026),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b26/B0_0 ));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_0_1  (
    .i0(inst_dob_i2_026),
    .i1(inst_dob_i3_026),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b26/B0_1 ));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_0_2  (
    .i0(inst_dob_i4_026),
    .i1(inst_dob_i5_026),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b26/B0_2 ));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_0_3  (
    .i0(inst_dob_i6_026),
    .i1(inst_dob_i7_026),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b26/B0_3 ));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b26/B0_0 ),
    .i1(\inst_dob_mux_b26/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b26/B1_0 ));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b26/B0_2 ),
    .i1(\inst_dob_mux_b26/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b26/B1_1 ));
  AL_MUX \inst_dob_mux_b26/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b26/B1_0 ),
    .i1(\inst_dob_mux_b26/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[26]));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_0_0  (
    .i0(inst_dob_i0_027),
    .i1(inst_dob_i0_027),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b27/B0_0 ));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_0_1  (
    .i0(inst_dob_i0_027),
    .i1(inst_dob_i0_027),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b27/B0_1 ));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_0_2  (
    .i0(inst_dob_i0_027),
    .i1(inst_dob_i0_027),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b27/B0_2 ));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_0_3  (
    .i0(inst_dob_i0_027),
    .i1(inst_dob_i0_027),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b27/B0_3 ));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b27/B0_0 ),
    .i1(\inst_dob_mux_b27/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b27/B1_0 ));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b27/B0_2 ),
    .i1(\inst_dob_mux_b27/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b27/B1_1 ));
  AL_MUX \inst_dob_mux_b27/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b27/B1_0 ),
    .i1(\inst_dob_mux_b27/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[27]));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_0_0  (
    .i0(inst_dob_i0_028),
    .i1(inst_dob_i0_028),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b28/B0_0 ));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_0_1  (
    .i0(inst_dob_i0_028),
    .i1(inst_dob_i0_028),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b28/B0_1 ));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_0_2  (
    .i0(inst_dob_i0_028),
    .i1(inst_dob_i0_028),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b28/B0_2 ));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_0_3  (
    .i0(inst_dob_i0_028),
    .i1(inst_dob_i0_028),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b28/B0_3 ));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b28/B0_0 ),
    .i1(\inst_dob_mux_b28/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b28/B1_0 ));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b28/B0_2 ),
    .i1(\inst_dob_mux_b28/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b28/B1_1 ));
  AL_MUX \inst_dob_mux_b28/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b28/B1_0 ),
    .i1(\inst_dob_mux_b28/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[28]));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_0_0  (
    .i0(inst_dob_i0_029),
    .i1(inst_dob_i0_029),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b29/B0_0 ));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_0_1  (
    .i0(inst_dob_i0_029),
    .i1(inst_dob_i0_029),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b29/B0_1 ));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_0_2  (
    .i0(inst_dob_i0_029),
    .i1(inst_dob_i0_029),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b29/B0_2 ));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_0_3  (
    .i0(inst_dob_i0_029),
    .i1(inst_dob_i0_029),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b29/B0_3 ));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b29/B0_0 ),
    .i1(\inst_dob_mux_b29/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b29/B1_0 ));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b29/B0_2 ),
    .i1(\inst_dob_mux_b29/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b29/B1_1 ));
  AL_MUX \inst_dob_mux_b29/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b29/B1_0 ),
    .i1(\inst_dob_mux_b29/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[29]));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_0  (
    .i0(inst_dob_i0_003),
    .i1(inst_dob_i1_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_1  (
    .i0(inst_dob_i2_003),
    .i1(inst_dob_i3_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_2  (
    .i0(inst_dob_i4_003),
    .i1(inst_dob_i5_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_3  (
    .i0(inst_dob_i6_003),
    .i1(inst_dob_i7_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b3/B0_0 ),
    .i1(\inst_dob_mux_b3/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b3/B0_2 ),
    .i1(\inst_dob_mux_b3/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b3/B1_0 ),
    .i1(\inst_dob_mux_b3/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[3]));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_0_0  (
    .i0(inst_dob_i0_030),
    .i1(inst_dob_i0_030),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b30/B0_0 ));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_0_1  (
    .i0(inst_dob_i0_030),
    .i1(inst_dob_i0_030),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b30/B0_1 ));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_0_2  (
    .i0(inst_dob_i0_030),
    .i1(inst_dob_i0_030),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b30/B0_2 ));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_0_3  (
    .i0(inst_dob_i0_030),
    .i1(inst_dob_i0_030),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b30/B0_3 ));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b30/B0_0 ),
    .i1(\inst_dob_mux_b30/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b30/B1_0 ));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b30/B0_2 ),
    .i1(\inst_dob_mux_b30/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b30/B1_1 ));
  AL_MUX \inst_dob_mux_b30/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b30/B1_0 ),
    .i1(\inst_dob_mux_b30/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[30]));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_0_0  (
    .i0(inst_dob_i0_031),
    .i1(inst_dob_i0_031),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b31/B0_0 ));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_0_1  (
    .i0(inst_dob_i0_031),
    .i1(inst_dob_i0_031),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b31/B0_1 ));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_0_2  (
    .i0(inst_dob_i0_031),
    .i1(inst_dob_i0_031),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b31/B0_2 ));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_0_3  (
    .i0(inst_dob_i0_031),
    .i1(inst_dob_i0_031),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b31/B0_3 ));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b31/B0_0 ),
    .i1(\inst_dob_mux_b31/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b31/B1_0 ));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b31/B0_2 ),
    .i1(\inst_dob_mux_b31/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b31/B1_1 ));
  AL_MUX \inst_dob_mux_b31/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b31/B1_0 ),
    .i1(\inst_dob_mux_b31/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[31]));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_0  (
    .i0(inst_dob_i0_004),
    .i1(inst_dob_i1_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_1  (
    .i0(inst_dob_i2_004),
    .i1(inst_dob_i3_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_2  (
    .i0(inst_dob_i4_004),
    .i1(inst_dob_i5_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_3  (
    .i0(inst_dob_i6_004),
    .i1(inst_dob_i7_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b4/B0_0 ),
    .i1(\inst_dob_mux_b4/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b4/B0_2 ),
    .i1(\inst_dob_mux_b4/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b4/B1_0 ),
    .i1(\inst_dob_mux_b4/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[4]));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_0  (
    .i0(inst_dob_i0_005),
    .i1(inst_dob_i1_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_1  (
    .i0(inst_dob_i2_005),
    .i1(inst_dob_i3_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_2  (
    .i0(inst_dob_i4_005),
    .i1(inst_dob_i5_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_3  (
    .i0(inst_dob_i6_005),
    .i1(inst_dob_i7_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b5/B0_0 ),
    .i1(\inst_dob_mux_b5/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b5/B0_2 ),
    .i1(\inst_dob_mux_b5/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b5/B1_0 ),
    .i1(\inst_dob_mux_b5/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[5]));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_0  (
    .i0(inst_dob_i0_006),
    .i1(inst_dob_i1_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_1  (
    .i0(inst_dob_i2_006),
    .i1(inst_dob_i3_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_2  (
    .i0(inst_dob_i4_006),
    .i1(inst_dob_i5_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_3  (
    .i0(inst_dob_i6_006),
    .i1(inst_dob_i7_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b6/B0_0 ),
    .i1(\inst_dob_mux_b6/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b6/B0_2 ),
    .i1(\inst_dob_mux_b6/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b6/B1_0 ),
    .i1(\inst_dob_mux_b6/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[6]));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_0  (
    .i0(inst_dob_i0_007),
    .i1(inst_dob_i1_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_1  (
    .i0(inst_dob_i2_007),
    .i1(inst_dob_i3_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_2  (
    .i0(inst_dob_i4_007),
    .i1(inst_dob_i5_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_3  (
    .i0(inst_dob_i6_007),
    .i1(inst_dob_i7_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b7/B0_0 ),
    .i1(\inst_dob_mux_b7/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b7/B0_2 ),
    .i1(\inst_dob_mux_b7/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b7/B1_0 ),
    .i1(\inst_dob_mux_b7/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[7]));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_0  (
    .i0(inst_dob_i0_008),
    .i1(inst_dob_i1_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_1  (
    .i0(inst_dob_i2_008),
    .i1(inst_dob_i3_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_2  (
    .i0(inst_dob_i4_008),
    .i1(inst_dob_i5_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_3  (
    .i0(inst_dob_i6_008),
    .i1(inst_dob_i7_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b8/B0_0 ),
    .i1(\inst_dob_mux_b8/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b8/B0_2 ),
    .i1(\inst_dob_mux_b8/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b8/B1_0 ),
    .i1(\inst_dob_mux_b8/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[8]));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_0  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i1_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_1  (
    .i0(inst_dob_i2_009),
    .i1(inst_dob_i3_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_2  (
    .i0(inst_dob_i4_009),
    .i1(inst_dob_i5_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_3  (
    .i0(inst_dob_i6_009),
    .i1(inst_dob_i7_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b9/B0_0 ),
    .i1(\inst_dob_mux_b9/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b9/B0_2 ),
    .i1(\inst_dob_mux_b9/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b9/B1_0 ),
    .i1(\inst_dob_mux_b9/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[9]));

endmodule 

