// Verilog netlist created by TD v4.6.116866
// Sat Nov 15 12:59:23 2025

`timescale 1ns / 1ps
module sample_memory  // al_ip/sample_memory.v(14)
  (
  addra,
  addrb,
  cea,
  clka,
  clkb,
  dia,
  dob
  );

  input [11:0] addra;  // al_ip/sample_memory.v(23)
  input [11:0] addrb;  // al_ip/sample_memory.v(24)
  input cea;  // al_ip/sample_memory.v(25)
  input clka;  // al_ip/sample_memory.v(26)
  input clkb;  // al_ip/sample_memory.v(27)
  input [31:0] dia;  // al_ip/sample_memory.v(22)
  output [31:0] dob;  // al_ip/sample_memory.v(19)


  // address_offset=0;data_offset=0;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_000 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n7,open_n8,open_n9,dia[1],open_n10,open_n11,dia[0],open_n12,open_n13}),
    .dob({open_n38,open_n39,open_n40,open_n41,open_n42,open_n43,open_n44,dob[1:0]}));
  // address_offset=0;data_offset=2;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_002 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n52,open_n53,open_n54,dia[3],open_n55,open_n56,dia[2],open_n57,open_n58}),
    .dob({open_n83,open_n84,open_n85,open_n86,open_n87,open_n88,open_n89,dob[3:2]}));
  // address_offset=0;data_offset=4;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_004 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n97,open_n98,open_n99,dia[5],open_n100,open_n101,dia[4],open_n102,open_n103}),
    .dob({open_n128,open_n129,open_n130,open_n131,open_n132,open_n133,open_n134,dob[5:4]}));
  // address_offset=0;data_offset=6;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_006 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n142,open_n143,open_n144,dia[7],open_n145,open_n146,dia[6],open_n147,open_n148}),
    .dob({open_n173,open_n174,open_n175,open_n176,open_n177,open_n178,open_n179,dob[7:6]}));
  // address_offset=0;data_offset=8;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_008 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n187,open_n188,open_n189,dia[9],open_n190,open_n191,dia[8],open_n192,open_n193}),
    .dob({open_n218,open_n219,open_n220,open_n221,open_n222,open_n223,open_n224,dob[9:8]}));
  // address_offset=0;data_offset=10;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_010 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n232,open_n233,open_n234,dia[11],open_n235,open_n236,dia[10],open_n237,open_n238}),
    .dob({open_n263,open_n264,open_n265,open_n266,open_n267,open_n268,open_n269,dob[11:10]}));
  // address_offset=0;data_offset=12;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_012 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n277,open_n278,open_n279,dia[13],open_n280,open_n281,dia[12],open_n282,open_n283}),
    .dob({open_n308,open_n309,open_n310,open_n311,open_n312,open_n313,open_n314,dob[13:12]}));
  // address_offset=0;data_offset=14;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_014 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n322,open_n323,open_n324,dia[15],open_n325,open_n326,dia[14],open_n327,open_n328}),
    .dob({open_n353,open_n354,open_n355,open_n356,open_n357,open_n358,open_n359,dob[15:14]}));
  // address_offset=0;data_offset=16;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_016 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n367,open_n368,open_n369,dia[17],open_n370,open_n371,dia[16],open_n372,open_n373}),
    .dob({open_n398,open_n399,open_n400,open_n401,open_n402,open_n403,open_n404,dob[17:16]}));
  // address_offset=0;data_offset=18;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_018 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n412,open_n413,open_n414,dia[19],open_n415,open_n416,dia[18],open_n417,open_n418}),
    .dob({open_n443,open_n444,open_n445,open_n446,open_n447,open_n448,open_n449,dob[19:18]}));
  // address_offset=0;data_offset=20;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_020 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n457,open_n458,open_n459,dia[21],open_n460,open_n461,dia[20],open_n462,open_n463}),
    .dob({open_n488,open_n489,open_n490,open_n491,open_n492,open_n493,open_n494,dob[21:20]}));
  // address_offset=0;data_offset=22;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_022 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n502,open_n503,open_n504,dia[23],open_n505,open_n506,dia[22],open_n507,open_n508}),
    .dob({open_n533,open_n534,open_n535,open_n536,open_n537,open_n538,open_n539,dob[23:22]}));
  // address_offset=0;data_offset=24;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_024 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n547,open_n548,open_n549,dia[25],open_n550,open_n551,dia[24],open_n552,open_n553}),
    .dob({open_n578,open_n579,open_n580,open_n581,open_n582,open_n583,open_n584,dob[25:24]}));
  // address_offset=0;data_offset=26;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_026 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n592,open_n593,open_n594,dia[27],open_n595,open_n596,dia[26],open_n597,open_n598}),
    .dob({open_n623,open_n624,open_n625,open_n626,open_n627,open_n628,open_n629,dob[27:26]}));
  // address_offset=0;data_offset=28;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_028 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n637,open_n638,open_n639,dia[29],open_n640,open_n641,dia[28],open_n642,open_n643}),
    .dob({open_n668,open_n669,open_n670,open_n671,open_n672,open_n673,open_n674,dob[29:28]}));
  // address_offset=0;data_offset=30;depth=4096;width=2;num_section=1;width_per_section=2;section_size=32;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x32_sub_000000_030 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .cea(cea),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n682,open_n683,open_n684,dia[31],open_n685,open_n686,dia[30],open_n687,open_n688}),
    .dob({open_n713,open_n714,open_n715,open_n716,open_n717,open_n718,open_n719,dob[31:30]}));

endmodule 

